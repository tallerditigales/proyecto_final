package arm_const;
	parameter VGA_SCREEN_SIZE = 160;
	parameter BLUE = 24'h0096FF;
	parameter WHITE = 24'hFFFFFF;
	parameter ORANGE = 24'hFD8000;
	parameter YELLOW = 24'hD1F523;
	parameter DARK = 24'h000000;
	parameter GREEN = 24'h228B22;
endpackage