package alu_defs;
//--------------------------------------------------------------------
// ALU RESULT TYPES
//--------------------------------------------------------------------
	parameter MOV_A =     2'b10;
	parameter MOV_B =     2'b11;
//--------------------------------------------------------------------
// ARITH_UNIT Operations
//--------------------------------------------------------------------
	parameter ARITH_ADD =  1'b0;
	parameter ARITH_SUB =  1'b1;
endpackage