module CPU_SINGLE_CYLCLE 
(

	input clk,
	input rst,
	input [31:0] instruction
	


);



endmodule