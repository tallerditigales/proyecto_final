package alu_defs;
//--------------------------------------------------------------------
// ALU RESULT TYPES
//--------------------------------------------------------------------
	parameter AND_ =     2'b10;
	parameter OR_ =     2'b11;
//--------------------------------------------------------------------
// ARITH_UNIT Operations
//--------------------------------------------------------------------
	parameter ARITH_ADD =  2'b00;
	parameter ARITH_SUB =  2'b01;
endpackage