module controller
(
	input logic clk, reset,
	input logic [31:12] Instr,
	input logic [3:0] ALUFlags,
	output logic [1:0] RegSrc,
	output logic RegWrite,
	output logic [1:0] ImmSrc,
	output logic ALUSrc,
	output logic [2:0] ALUControl,
	output logic MemWrite, MemtoReg,
	output logic PCSrc
);

	logic [1:0] FlagW;
	logic PCS, RegW, MemW;
	
	// MEMORY	
	// 								   	 FUNCT																	 11:0
	//	31:28	  27:26	  	-------------25:20-------------	 19:16  	 15:12   	  11:0	 ->	imm12 
	//	cond		op			I		P		U		B		W		L		Rn			Rd				Src	 		
	//																												 ->	shamt5|sh| 1 |Rm
	//																														 11:7	 6:5 4  3:0
	
	decoder dec(Instr[27:26], Instr[25:20], Instr[15:12],
					FlagW, PCS, RegW, MemW,
					MemtoReg, ALUSrc, ImmSrc, 
					RegSrc, ALUControl);
	
	condlogic cl(clk, reset, Instr[31:28], ALUFlags,
					FlagW, PCS, RegW, MemW,
					PCSrc, RegWrite, MemWrite);
					
endmodule